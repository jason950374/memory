sram_8T

.subckt sram_8T WWL RWL WBL WBL_B RBL nVdd
Mp_inv1 		nData	nData_b	nVdd	nVdd
Mp_inv2 		nData_b	nData	nVdd	nVdd
Mn_inv1 		nData	nData_b	gnd		gnd
Mn_inv2 		nData_b	nData	gnd		gnd
Mn_W_PG			nData	WWL		WBL		gnd
Mn_W_PG_b		nData_b	WWL		WBL_B	gnd
Mn_R_PullDown	nTemp	nData	gnd		gnd
Mn_R_PG			RBL		RWL		nTemp		gnd
.ends

















